# ====================================================================
#
#      audio_arm_dadio.cdl
#
#      eCos audio layer for iobjects dadio
#
# ====================================================================
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      toddm
# Original data:  toddm
# Contributors:   ericg danb
# Date:           2000-12-09
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package DDOPKG_IO_AUDIO_ARM_DADIO {
    display       "Dadio Maverick Audio - CS4341 DAC"
#    parent	  DDOPKG_IO_AUDIO_ARM_DADIO
    include_dir	  dadio/io
    include_files audio.h audio_asm.h i2c.h
    description   "
        This option enables the driver for Dadio players based on Cirrus Logic's Maverick
      	part."
#    doc           redirect/ecos-device-drivers.html

    compile       -library=libextras.a   audio.c i2c.c i2s_fiq.S

    cdl_option DDODAT_IO_AUDIO_NAME {
	display		"Audio device name"
	flavor		data
	default_value	{ "\"/dev/dsp\"" }
	description	"
	    The name of the Audio device."
    } 

    cdl_component DDOPKG_IO_AUDIO_ARM_DADIO_OPTIONS {
        display "Audio build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option DDOPKG_IO_AUDIO_ARM_DADIO_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option DDOPKG_IO_AUDIO_ARM_DADIO_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }

	cdl_option DDOPKG_IO_AUDIO_ARM_DADIO_TESTS {
	    display "Audio tests"
 	    flavor  data
            no_define
            calculated { "tests/audio_test" }
	    description "
                This option specifies the set of tests for the Audio HW."
	}
    }
}

# EOF audio_arm_dadio.cdl



