# ====================================================================
#
#      usb_arm_dadio.cdl
#
#      eCos usb layer for iobjects dadio
#
# ====================================================================
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      toddm
# Original data:  toddm
# Contributors:
# Date:           2000-07-26
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package DDOPKG_IO_USB_ARM_DADIO {
    display       "Dadio USB driver"
#    parent	  DDOPKG_DADIO
    include_dir	  dadio/io
    include_files usb.h
    description   "
        This option enables the usb driver."
#    doc           redirect/ecos-device-drivers.html

    compile       -library=libextras.a   usb.c

    cdl_option DDODAT_IO_USB_NAME {
	display		"USB device name"
	flavor		data
	default_value	{ "\"/dev/usb\"" }
	description	"
		This option includes the USB driver for the Mystic chip."
    }

    cdl_component DDOPKG_IO_USB_ARM_DADIO_OPTIONS {
        display "USB build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option DDOPKG_IO_USB_ARM_DADIO_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are used in addition
                to the set of global flags."
        }

        cdl_option DDOPKG_IO_USB_ARM_DADIO_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building these serial device drivers. These flags are removed from
                the set of global flags if present."
        }

	cdl_option DDOPKG_IO_USB_ARM_DADIO_TESTS {
	    display "USB tests"
 	    flavor  data
            no_define
            calculated { "tests/usb_test" }
	    description "
                This option specifies the set of tests for the USB
               driver."
	}
    }
}

# EOF usb_arm_dadio.cdl



