# ====================================================================
#
#      lcd_arm_dadio.cdl
#
#      eCos lcd layer for iobjects dadio
#
# ====================================================================
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      toddm
# Original data:  toddm
# Contributors:
# Date:           2000-06-09
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package DDOPKG_IO_LCD_ARM_DADIO {
    display       "Dadio LCD driver"
#    parent	  DDOPKG_DADIO
    include_dir	  dadio/io
    include_files lcd.h
    description   "
        This option enables the power management sub-system."
#    doc           redirect/ecos-device-drivers.html

    compile       -library=libextras.a   lcd.c

    cdl_option DDODAT_IO_LCD_NAME {
	display		"LCD device name"
	flavor		data
	default_value	{ "\"/dev/lcd\"" }
	description	"
		Getting a handle to this device allows access to the LCD."
    }

    cdl_component DDOPKG_IO_LCD_ARM_DADIO_OPTIONS {
        display "LCD build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option DDOPKG_IO_LCD_ARM_DADIO_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this LCD driver. These flags are used in addition
                to the set of global flags."
        }

        cdl_option DDOPKG_IO_LCD_ARM_DADIO_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building this LCD driver. These flags are removed from
                the set of global flags if present."
        }

	cdl_option DDOPKG_IO_LCD_ARM_DADIO_TESTS {
	    display "LCD tests"
 	    flavor  data
            no_define
            calculated { "tests/lcd_test" }
	    description "
                This option specifies the set of tests for the LCD driver."
	}
    }
}

# EOF lcd_arm_dadio.cdl
